interface ClkDivBy2;
logic en,clk,rst;
logic div2,div4,div8,div16;
endinterface