interface A_C ;
logic [3:0] A,B;
logic m;
logic [4:0] result;
endinterface