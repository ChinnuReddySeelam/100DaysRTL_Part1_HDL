module FA(input a, b, cin, output sum, carry);  assign {carry, sum} = a + b + cin;endmodulemodule A_S(  input [3:0] A, B,  input m,  output [4:0] result,  output overflow);wire [3:0] Y;wire [3:0] C;wire [3:0] S;wire cout_sub;xor X1(Y[0],m,B[0]);xor X2(Y[1],m,B[1]);xor X3(Y[2],m,B[2]);xor X4(Y[3],m,B[3]);FA FA1(A[0], Y[0], m, S[0], C[0]);FA FA2(A[1], Y[1], C[0], S[1], C[1]);FA FA3(A[2], Y[2], C[1], S[2], C[2]);FA FA4(A[3], Y[3], C[2], S[3], C[3]);assign overflow = ((A[3] & Y[3] & ~S[3]) | (~A[3] & ~Y[3] & S[3])) | cout_sub;assign cout_sub = (m == 1'b1) ? ~C[3] : C[3];assign result = {cout_sub, S};endmodule