interface Clk_Div_by_odd;
logic clk,rst;
logic div3,div5,div9;
endinterface